library verilog;
use verilog.vl_types.all;
entity somethingIsWrong is
    port(
        somethingiswrong: out    vl_logic;
        bigbombpossible : in     vl_logic;
        validlocation   : in     vl_logic
    );
end somethingIsWrong;
