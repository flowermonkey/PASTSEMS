library verilog;
use verilog.vl_types.all;
entity Battleship_sv_unit is
end Battleship_sv_unit;
