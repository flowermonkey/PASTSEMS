library verilog;
use verilog.vl_types.all;
entity BCDtoSevenSeg is
    port(
        led             : out    vl_logic_vector(7 downto 0);
        bcd             : in     vl_logic_vector(3 downto 0)
    );
end BCDtoSevenSeg;
