library verilog;
use verilog.vl_types.all;
entity library_sv_unit is
end library_sv_unit;
