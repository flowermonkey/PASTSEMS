
module priQueue ( newVal, ck, r, clear, loadIn, shiftOut, top );
  input [7:0] newVal;
  output [7:0] top;
  input ck, r, clear, loadIn, shiftOut;
  wire   \r6/N1 , n14, n17, n20, n23, n26, n29, n32, n35, n38, n41, n44, n47,
         n50, n53, n56, n59, n62, n65, n68, n71, n74, n77, n80, n83, n86, n89,
         n92, n95, n98, n101, n104, n107, n110, n113, n116, n119, n122, n125,
         n128, n131, n134, n137, n140, n143, n146, n149, n152, n156, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n918,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n935, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n951, n952, n953, n954, n955, n956,
         n957, n960, n961, n962, n963, n964, n966, n967, n968, n969, n970,
         n971, n972, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n987, n988, n989, n990, n991, n993, n994, n995, n996,
         n997, n998, n1000, n1001, n1002, n1003, n1004, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1030, n1031, n1039, n1045,
         n1046, n1047, n1048, n1049, n1050, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1063, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1075, n1076, n1077, n1078, n1079,
         n1080, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168;
  wire   [7:0] r2_out;
  wire   [7:0] r3_out;
  wire   [7:0] r4_out;
  wire   [7:0] r5_out;
  wire   [7:0] r6_out;
  assign \r6/N1  = r;

  DFFSX1 \r5/out_reg[7]  ( .D(n128), .CK(ck), .SN(n1168), .Q(n1166), .QN(
        r5_out[7]) );
  DFFSX1 \r3/out_reg[7]  ( .D(n122), .CK(ck), .SN(n1168), .Q(n1165), .QN(
        r3_out[7]) );
  DFFSX1 \r6/out_reg[4]  ( .D(n62), .CK(ck), .SN(n1168), .Q(n1164), .QN(
        r6_out[4]) );
  DFFSX1 \r3/out_reg[2]  ( .D(n32), .CK(ck), .SN(n1168), .Q(n1163), .QN(
        r3_out[2]) );
  DFFSX1 \r4/out_reg[5]  ( .D(n86), .CK(ck), .SN(n1168), .Q(n1162), .QN(
        r4_out[5]) );
  DFFSX1 \r1/out_reg[6]  ( .D(n89), .CK(ck), .SN(n1168), .Q(n1161), .QN(top[6]) );
  DFFSX1 \r4/out_reg[4]  ( .D(n68), .CK(ck), .SN(n1168), .Q(n1160), .QN(
        r4_out[4]) );
  DFFSX1 \r5/out_reg[3]  ( .D(n47), .CK(ck), .SN(n1168), .Q(n1159), .QN(
        r5_out[3]) );
  DFFSX1 \r4/out_reg[3]  ( .D(n50), .CK(ck), .SN(n1168), .Q(n1158), .QN(
        r4_out[3]) );
  DFFSX1 \r3/out_reg[6]  ( .D(n95), .CK(ck), .SN(n1168), .Q(n1157), .QN(
        r3_out[6]) );
  DFFSX1 \r1/out_reg[7]  ( .D(n152), .CK(ck), .SN(n1168), .Q(n1156), .QN(
        top[7]) );
  DFFSX1 \r2/out_reg[5]  ( .D(n74), .CK(ck), .SN(n1168), .Q(n1155), .QN(
        r2_out[5]) );
  DFFSX1 \r1/out_reg[2]  ( .D(n110), .CK(ck), .SN(n1168), .Q(n1154), .QN(
        top[2]) );
  DFFSX1 \r2/out_reg[3]  ( .D(n38), .CK(ck), .SN(n1168), .Q(n1153), .QN(
        r2_out[3]) );
  DFFSX1 \r6/out_reg[6]  ( .D(n98), .CK(ck), .SN(n1168), .QN(r6_out[6]) );
  DFFSX1 \r6/out_reg[5]  ( .D(n80), .CK(ck), .SN(n1168), .QN(r6_out[5]) );
  DFFSX1 \r6/out_reg[7]  ( .D(n131), .CK(ck), .SN(n1168), .QN(r6_out[7]) );
  DFFSX1 \r5/out_reg[6]  ( .D(n101), .CK(ck), .SN(n1168), .QN(r5_out[6]) );
  DFFSX1 \r6/out_reg[1]  ( .D(n17), .CK(ck), .SN(n1168), .QN(r6_out[1]) );
  DFFSX1 \r1/out_reg[4]  ( .D(n53), .CK(ck), .SN(n1168), .QN(top[4]) );
  DFFSX1 \r6/out_reg[2]  ( .D(n23), .CK(ck), .SN(n1168), .QN(r6_out[2]) );
  DFFSX1 \r3/out_reg[1]  ( .D(n116), .CK(ck), .SN(n1168), .QN(r3_out[1]) );
  DFFSX1 \r5/out_reg[2]  ( .D(n26), .CK(ck), .SN(n1168), .QN(r5_out[2]) );
  DFFSX1 \r2/out_reg[6]  ( .D(n92), .CK(ck), .SN(n1168), .QN(r2_out[6]) );
  DFFSX1 \r2/out_reg[7]  ( .D(n156), .CK(ck), .SN(n1168), .QN(r2_out[7]) );
  DFFSX1 \r4/out_reg[2]  ( .D(n29), .CK(ck), .SN(n1168), .QN(r4_out[2]) );
  DFFSX1 \r3/out_reg[0]  ( .D(n143), .CK(ck), .SN(n1168), .QN(r3_out[0]) );
  DFFSX1 \r5/out_reg[1]  ( .D(n20), .CK(ck), .SN(n1168), .QN(r5_out[1]) );
  DFFSX1 \r4/out_reg[1]  ( .D(n113), .CK(ck), .SN(n1168), .QN(r4_out[1]) );
  DFFSX1 \r3/out_reg[4]  ( .D(n59), .CK(ck), .SN(n1168), .QN(r3_out[4]) );
  DFFSX1 \r1/out_reg[5]  ( .D(n71), .CK(ck), .SN(n1168), .QN(top[5]) );
  DFFSX1 \r6/out_reg[0]  ( .D(n134), .CK(ck), .SN(n1168), .QN(r6_out[0]) );
  DFFSX1 \r5/out_reg[5]  ( .D(n83), .CK(ck), .SN(n1168), .QN(r5_out[5]) );
  DFFSX1 \r2/out_reg[4]  ( .D(n56), .CK(ck), .SN(n1168), .QN(r2_out[4]) );
  DFFSX1 \r6/out_reg[3]  ( .D(n44), .CK(ck), .SN(n1168), .QN(r6_out[3]) );
  DFFSX1 \r5/out_reg[4]  ( .D(n65), .CK(ck), .SN(n1168), .QN(r5_out[4]) );
  DFFSX1 \r4/out_reg[6]  ( .D(n104), .CK(ck), .SN(n1168), .QN(r4_out[6]) );
  DFFSX1 \r4/out_reg[0]  ( .D(n140), .CK(ck), .SN(n1168), .QN(r4_out[0]) );
  DFFSX1 \r4/out_reg[7]  ( .D(n125), .CK(ck), .SN(n1168), .QN(r4_out[7]) );
  DFFSX1 \r3/out_reg[5]  ( .D(n77), .CK(ck), .SN(n1168), .QN(r3_out[5]) );
  DFFSX1 \r5/out_reg[0]  ( .D(n137), .CK(ck), .SN(n1168), .QN(r5_out[0]) );
  DFFSX1 \r3/out_reg[3]  ( .D(n41), .CK(ck), .SN(n1168), .QN(r3_out[3]) );
  DFFSX1 \r1/out_reg[1]  ( .D(n14), .CK(ck), .SN(n1168), .QN(top[1]) );
  DFFSX1 \r1/out_reg[0]  ( .D(n149), .CK(ck), .SN(n1168), .QN(top[0]) );
  DFFSX1 \r2/out_reg[2]  ( .D(n107), .CK(ck), .SN(n1168), .QN(r2_out[2]) );
  DFFSX1 \r2/out_reg[1]  ( .D(n119), .CK(ck), .SN(n1168), .QN(r2_out[1]) );
  DFFSX1 \r1/out_reg[3]  ( .D(n35), .CK(ck), .SN(n1168), .QN(top[3]) );
  DFFSX1 \r2/out_reg[0]  ( .D(n146), .CK(ck), .SN(n1168), .QN(r2_out[0]) );
  OAI21XL U734 ( .A0(r2_out[0]), .A1(n1012), .B0(r2_out[1]), .Y(n1084) );
  OAI21XL U639 ( .A0(r6_out[0]), .A1(n1012), .B0(r6_out[1]), .Y(n1010) );
  OAI21XL U636 ( .A0(r6_out[3]), .A1(n951), .B0(n1007), .Y(n1006) );
  OAI222XL U633 ( .A0(n1003), .A1(n1004), .B0(r6_out[6]), .B1(n920), .C0(
        r6_out[5]), .C1(n937), .Y(n1002) );
  OAI22XL U701 ( .A0(r4_out[7]), .A1(n960), .B0(r4_out[6]), .B1(n920), .Y(
        n1048) );
  AOI211XL U699 ( .A0(r4_out[3]), .A1(n951), .B0(r4_out[2]), .C0(n987), .Y(
        n1054) );
  OAI21XL U696 ( .A0(r4_out[0]), .A1(n1012), .B0(r4_out[1]), .Y(n1058) );
  OAI21XL U695 ( .A0(n1158), .A1(newVal[3]), .B0(n1058), .Y(n1057) );
  AOI211XL U694 ( .A0(r4_out[2]), .A1(n987), .B0(n1056), .C0(n1057), .Y(n1055)
         );
  OAI21XL U692 ( .A0(r4_out[3]), .A1(n951), .B0(n1053), .Y(n1052) );
  NOR3X1 U583 ( .A(n967), .B(n969), .C(n966), .Y(n906) );
  AOI2BB2XL U577 ( .B0(r5_out[0]), .B1(n929), .A0N(n964), .A1N(n910), .Y(n137)
         );
  AOI2BB2XL U526 ( .B0(r5_out[5]), .B1(n929), .A0N(n930), .A1N(n910), .Y(n83)
         );
  AOI2BB2XL U547 ( .B0(r5_out[3]), .B1(n929), .A0N(n947), .A1N(n910), .Y(n47)
         );
  AOI2BB2XL U560 ( .B0(r5_out[2]), .B1(n929), .A0N(n955), .A1N(n910), .Y(n26)
         );
  AOI222XL U588 ( .A0(n931), .A1(r4_out[7]), .B0(n911), .B1(r6_out[7]), .C0(
        newVal[7]), .C1(n932), .Y(n974) );
  AOI2BB2XL U587 ( .B0(r5_out[7]), .B1(n929), .A0N(n974), .A1N(n910), .Y(n128)
         );
  AOI2BB2XL U537 ( .B0(r5_out[4]), .B1(n929), .A0N(n943), .A1N(n910), .Y(n65)
         );
  AOI2BB2XL U563 ( .B0(r5_out[1]), .B1(n929), .A0N(n956), .A1N(n910), .Y(n20)
         );
  AOI222XL U623 ( .A0(n931), .A1(r4_out[6]), .B0(n911), .B1(r6_out[6]), .C0(
        newVal[6]), .C1(n932), .Y(n994) );
  AOI2BB2XL U622 ( .B0(r5_out[6]), .B1(n929), .A0N(n994), .A1N(n910), .Y(n101)
         );
  OAI222XL U607 ( .A0(loadIn), .A1(n1163), .B0(n918), .B1(n1154), .C0(n987), 
        .C1(n921), .Y(n984) );
  OAI222XL U522 ( .A0(loadIn), .A1(n1157), .B0(n918), .B1(n1161), .C0(n920), 
        .C1(n921), .Y(n915) );
  AOI22XL U521 ( .A0(r2_out[6]), .A1(n914), .B0(n915), .B1(n1167), .Y(n92) );
  OAI222XL U567 ( .A0(loadIn), .A1(n1165), .B0(n918), .B1(n1156), .C0(n960), 
        .C1(n921), .Y(n957) );
  AOI22XL U566 ( .A0(r2_out[7]), .A1(n914), .B0(n957), .B1(n1167), .Y(n156) );
  AOI2BB2XL U570 ( .B0(r2_out[0]), .B1(n914), .A0N(n961), .A1N(n910), .Y(n146)
         );
  AOI2BB2XL U593 ( .B0(r2_out[1]), .B1(n914), .A0N(n977), .A1N(n910), .Y(n119)
         );
  AOI2BB2XL U542 ( .B0(r2_out[4]), .B1(n914), .A0N(n945), .A1N(n910), .Y(n56)
         );
  AOI2BB2XL U532 ( .B0(r2_out[5]), .B1(n914), .A0N(n939), .A1N(n910), .Y(n74)
         );
  AOI2BB2XL U553 ( .B0(r2_out[3]), .B1(n914), .A0N(n952), .A1N(n910), .Y(n38)
         );
  AOI222XL U590 ( .A0(n927), .A1(r3_out[7]), .B0(n911), .B1(r5_out[7]), .C0(
        newVal[7]), .C1(n928), .Y(n975) );
  AOI2BB2XL U589 ( .B0(r4_out[7]), .B1(n925), .A0N(n975), .A1N(n910), .Y(n125)
         );
  AOI222XL U575 ( .A0(n927), .A1(r3_out[0]), .B0(n911), .B1(r5_out[0]), .C0(
        newVal[0]), .C1(n928), .Y(n963) );
  AOI2BB2XL U574 ( .B0(r4_out[0]), .B1(n925), .A0N(n963), .A1N(n910), .Y(n140)
         );
  AOI222XL U612 ( .A0(n927), .A1(r3_out[6]), .B0(n911), .B1(r5_out[6]), .C0(
        newVal[6]), .C1(n928), .Y(n988) );
  AOI2BB2XL U611 ( .B0(r4_out[6]), .B1(n925), .A0N(n988), .A1N(n910), .Y(n104)
         );
  AOI222XL U546 ( .A0(n927), .A1(r3_out[3]), .B0(n911), .B1(r5_out[3]), .C0(
        newVal[3]), .C1(n928), .Y(n946) );
  AOI2BB2XL U545 ( .B0(r4_out[3]), .B1(n925), .A0N(n946), .A1N(n910), .Y(n50)
         );
  AOI222XL U601 ( .A0(n927), .A1(r3_out[1]), .B0(n911), .B1(r5_out[1]), .C0(
        newVal[1]), .C1(n928), .Y(n982) );
  AOI2BB2XL U600 ( .B0(r4_out[1]), .B1(n925), .A0N(n982), .A1N(n910), .Y(n113)
         );
  AOI222XL U525 ( .A0(n927), .A1(r3_out[5]), .B0(n911), .B1(r5_out[5]), .C0(
        newVal[5]), .C1(n928), .Y(n926) );
  AOI2BB2XL U524 ( .B0(r4_out[5]), .B1(n925), .A0N(n926), .A1N(n910), .Y(n86)
         );
  AOI222XL U559 ( .A0(n927), .A1(r3_out[2]), .B0(n911), .B1(r5_out[2]), .C0(
        newVal[2]), .C1(n928), .Y(n954) );
  AOI2BB2XL U558 ( .B0(r4_out[2]), .B1(n925), .A0N(n954), .A1N(n910), .Y(n29)
         );
  AOI222XL U536 ( .A0(n927), .A1(r3_out[4]), .B0(n911), .B1(r5_out[4]), .C0(
        newVal[4]), .C1(n928), .Y(n942) );
  AOI2BB2XL U535 ( .B0(r4_out[4]), .B1(n925), .A0N(n942), .A1N(n910), .Y(n68)
         );
  OAI222XL U551 ( .A0(loadIn), .A1(n1158), .B0(n935), .B1(n1153), .C0(n951), 
        .C1(n938), .Y(n948) );
  OAI222XL U531 ( .A0(loadIn), .A1(n1162), .B0(n935), .B1(n1155), .C0(n937), 
        .C1(n938), .Y(n933) );
  AOI222XL U592 ( .A0(n911), .A1(r4_out[7]), .B0(n912), .B1(r2_out[7]), .C0(
        newVal[7]), .C1(n913), .Y(n976) );
  AOI2BB2XL U591 ( .B0(r3_out[7]), .B1(n908), .A0N(n976), .A1N(n910), .Y(n122)
         );
  AOI222XL U573 ( .A0(n911), .A1(r4_out[0]), .B0(n912), .B1(r2_out[0]), .C0(
        newVal[0]), .C1(n913), .Y(n962) );
  AOI2BB2XL U572 ( .B0(r3_out[0]), .B1(n908), .A0N(n962), .A1N(n910), .Y(n143)
         );
  AOI222XL U557 ( .A0(n911), .A1(r4_out[2]), .B0(n912), .B1(r2_out[2]), .C0(
        newVal[2]), .C1(n913), .Y(n953) );
  AOI2BB2XL U556 ( .B0(r3_out[2]), .B1(n908), .A0N(n953), .A1N(n910), .Y(n32)
         );
  AOI222XL U520 ( .A0(n911), .A1(r4_out[6]), .B0(n912), .B1(r2_out[6]), .C0(
        newVal[6]), .C1(n913), .Y(n909) );
  AOI2BB2XL U519 ( .B0(r3_out[6]), .B1(n908), .A0N(n909), .A1N(n910), .Y(n95)
         );
  AOI222XL U597 ( .A0(n911), .A1(r4_out[1]), .B0(n912), .B1(r2_out[1]), .C0(
        newVal[1]), .C1(n913), .Y(n978) );
  AOI2BB2XL U596 ( .B0(r3_out[1]), .B1(n908), .A0N(n978), .A1N(n910), .Y(n116)
         );
  AOI222XL U541 ( .A0(n911), .A1(r4_out[4]), .B0(n912), .B1(r2_out[4]), .C0(
        newVal[4]), .C1(n913), .Y(n944) );
  AOI2BB2XL U540 ( .B0(r3_out[4]), .B1(n908), .A0N(n944), .A1N(n910), .Y(n59)
         );
  AOI222XL U523 ( .A0(n922), .A1(top[6]), .B0(r2_out[6]), .B1(n923), .C0(
        newVal[6]), .C1(n924), .Y(n89) );
  AOI222XL U568 ( .A0(n922), .A1(top[7]), .B0(r2_out[7]), .B1(n923), .C0(
        newVal[7]), .C1(n924), .Y(n152) );
  NAND2X1 U614 ( .A(loadIn), .B(n991), .Y(n980) );
  NAND2X1 U743 ( .A(newVal[5]), .B(n1155), .Y(n1076) );
  OAI211X1 U733 ( .A0(n1082), .A1(newVal[1]), .B0(n1083), .C0(n1084), .Y(n1080) );
  AOI211X1 U729 ( .A0(newVal[3]), .A1(n1153), .B0(n1078), .C0(n1079), .Y(n1077) );
  AOI222X1 U635 ( .A0(newVal[4]), .A1(n1164), .B0(n1164), .B1(n1006), .C0(
        newVal[4]), .C1(n1006), .Y(n1003) );
  AOI2BB1XL U719 ( .A0N(n1013), .A1N(top[0]), .B0(newVal[1]), .Y(n1070) );
  AOI211X1 U717 ( .A0(top[1]), .A1(n1069), .B0(n1070), .C0(n1071), .Y(n1067)
         );
  AOI222X1 U714 ( .A0(n1067), .A1(n1154), .B0(n1067), .B1(newVal[2]), .C0(
        n1154), .C1(n1068), .Y(n1066) );
  AOI2BB1XL U711 ( .A0N(newVal[4]), .A1N(n1063), .B0(top[4]), .Y(n1065) );
  AOI2BB1XL U698 ( .A0N(n1013), .A1N(r4_out[0]), .B0(newVal[1]), .Y(n1056) );
  AOI2BB1XL U688 ( .A0N(r4_out[7]), .A1N(n1045), .B0(newVal[7]), .Y(n1047) );
  NOR3X1 U629 ( .A(n997), .B(n967), .C(n998), .Y(n970) );
  INVX1 U621 ( .A(n981), .Y(n968) );
  NAND2X1 U628 ( .A(loadIn), .B(n996), .Y(n995) );
  NOR2X1 U609 ( .A(n983), .B(n935), .Y(n941) );
  INVX1 U608 ( .A(n941), .Y(n921) );
  NOR3X1 U613 ( .A(n989), .B(n990), .C(n980), .Y(n928) );
  INVX1 U552 ( .A(n913), .Y(n938) );
  NAND2X1 U646 ( .A(loadIn), .B(n1167), .Y(n969) );
  AOI222XL U518 ( .A0(n905), .A1(r5_out[6]), .B0(newVal[6]), .B1(n906), .C0(
        n907), .C1(r6_out[6]), .Y(n98) );
  AOI222XL U579 ( .A0(n905), .A1(r5_out[0]), .B0(newVal[0]), .B1(n906), .C0(
        n907), .C1(r6_out[0]), .Y(n134) );
  AOI222XL U529 ( .A0(n905), .A1(r5_out[5]), .B0(newVal[5]), .B1(n906), .C0(
        n907), .C1(r6_out[5]), .Y(n80) );
  AOI222XL U580 ( .A0(n905), .A1(r5_out[7]), .B0(newVal[7]), .B1(n906), .C0(
        n907), .C1(r6_out[7]), .Y(n131) );
  AOI222XL U539 ( .A0(n905), .A1(r5_out[4]), .B0(newVal[4]), .B1(n906), .C0(
        n907), .C1(r6_out[4]), .Y(n62) );
  AOI222XL U565 ( .A0(n905), .A1(r5_out[1]), .B0(newVal[1]), .B1(n906), .C0(
        n907), .C1(r6_out[1]), .Y(n17) );
  AOI222XL U562 ( .A0(n905), .A1(r5_out[2]), .B0(newVal[2]), .B1(n906), .C0(
        n907), .C1(r6_out[2]), .Y(n23) );
  AOI222XL U549 ( .A0(n905), .A1(r5_out[3]), .B0(newVal[3]), .B1(n906), .C0(
        n907), .C1(r6_out[3]), .Y(n44) );
  AOI222XL U578 ( .A0(n931), .A1(r4_out[0]), .B0(n911), .B1(r6_out[0]), .C0(
        newVal[0]), .C1(n932), .Y(n964) );
  AOI222XL U527 ( .A0(n931), .A1(r4_out[5]), .B0(n911), .B1(r6_out[5]), .C0(
        newVal[5]), .C1(n932), .Y(n930) );
  AOI222XL U548 ( .A0(n931), .A1(r4_out[3]), .B0(n911), .B1(r6_out[3]), .C0(
        newVal[3]), .C1(n932), .Y(n947) );
  AOI222XL U561 ( .A0(n931), .A1(r4_out[2]), .B0(n911), .B1(r6_out[2]), .C0(
        newVal[2]), .C1(n932), .Y(n955) );
  AOI222XL U538 ( .A0(n931), .A1(r4_out[4]), .B0(n911), .B1(r6_out[4]), .C0(
        newVal[4]), .C1(n932), .Y(n943) );
  AOI222XL U564 ( .A0(n931), .A1(r4_out[1]), .B0(n911), .B1(r6_out[1]), .C0(
        newVal[1]), .C1(n932), .Y(n956) );
  AOI222XL U571 ( .A0(n911), .A1(r3_out[0]), .B0(n940), .B1(top[0]), .C0(
        newVal[0]), .C1(n941), .Y(n961) );
  AOI222XL U594 ( .A0(n911), .A1(r3_out[1]), .B0(n940), .B1(top[1]), .C0(
        newVal[1]), .C1(n941), .Y(n977) );
  AOI222XL U543 ( .A0(n911), .A1(r3_out[4]), .B0(n940), .B1(top[4]), .C0(
        newVal[4]), .C1(n941), .Y(n945) );
  AOI222XL U533 ( .A0(n911), .A1(r3_out[5]), .B0(n940), .B1(top[5]), .C0(
        newVal[5]), .C1(n941), .Y(n939) );
  AOI222XL U554 ( .A0(n911), .A1(r3_out[3]), .B0(n940), .B1(top[3]), .C0(
        newVal[3]), .C1(n941), .Y(n952) );
  AOI222XL U555 ( .A0(n922), .A1(top[3]), .B0(r2_out[3]), .B1(n923), .C0(
        newVal[3]), .C1(n924), .Y(n35) );
  AOI222XL U544 ( .A0(n922), .A1(top[4]), .B0(r2_out[4]), .B1(n923), .C0(
        newVal[4]), .C1(n924), .Y(n53) );
  AOI222XL U569 ( .A0(n922), .A1(top[0]), .B0(r2_out[0]), .B1(n923), .C0(
        newVal[0]), .C1(n924), .Y(n149) );
  AOI222XL U534 ( .A0(n922), .A1(top[5]), .B0(r2_out[5]), .B1(n923), .C0(
        newVal[5]), .C1(n924), .Y(n71) );
  AOI222XL U576 ( .A0(n922), .A1(top[1]), .B0(r2_out[1]), .B1(n923), .C0(
        newVal[1]), .C1(n924), .Y(n14) );
  AOI222XL U602 ( .A0(n922), .A1(top[2]), .B0(r2_out[2]), .B1(n923), .C0(
        newVal[2]), .C1(n924), .Y(n110) );
  AOI21XL U690 ( .A0(r4_out[5]), .A1(n937), .B0(n1050), .Y(n1049) );
  AOI211XL U687 ( .A0(r4_out[7]), .A1(n1045), .B0(n1046), .C0(n1047), .Y(n1031) );
  NOR2XL U740 ( .A(r2_out[4]), .B(n1030), .Y(n1078) );
  NOR2BX1 U718 ( .AN(top[3]), .B(newVal[3]), .Y(n1071) );
  AOI22XL U530 ( .A0(r3_out[5]), .A1(n908), .B0(n933), .B1(n1167), .Y(n77) );
  AOI21XL U715 ( .A0(top[3]), .A1(n951), .B0(n987), .Y(n1068) );
  NOR2BX1 U634 ( .AN(r6_out[5]), .B(newVal[5]), .Y(n1004) );
  AOI211XL U638 ( .A0(r6_out[3]), .A1(n951), .B0(r6_out[2]), .C0(n987), .Y(
        n1011) );
  OR2X1 U720 ( .A(n1012), .B(top[0]), .Y(n1069) );
  AOI22XL U640 ( .A0(r6_out[3]), .A1(n951), .B0(n1013), .B1(n1014), .Y(n1009)
         );
  AOI22XL U641 ( .A0(r6_out[0]), .A1(n1014), .B0(r6_out[2]), .B1(n987), .Y(
        n1008) );
  NOR2XL U738 ( .A(n1013), .B(r2_out[0]), .Y(n1082) );
  NAND2XL U736 ( .A(r2_out[3]), .B(n951), .Y(n1083) );
  AOI31XL U637 ( .A0(n1008), .A1(n1009), .A2(n1010), .B0(n1011), .Y(n1007) );
  AOI211XL U693 ( .A0(newVal[4]), .A1(n1160), .B0(n1054), .C0(n1055), .Y(n1053) );
  AOI32X1 U728 ( .A0(r2_out[4]), .A1(n1076), .A2(n1030), .B0(n1077), .B1(n1076), .Y(n1075) );
  OAI2BB1X1 U632 ( .A0N(r6_out[6]), .A1N(n920), .B0(n1002), .Y(n1001) );
  AOI211XL U689 ( .A0(newVal[5]), .A1(n1162), .B0(n1048), .C0(n1049), .Y(n1046) );
  OR2X2 U669 ( .A(n1031), .B(n989), .Y(n998) );
  AOI22XL U550 ( .A0(r3_out[3]), .A1(n908), .B0(n948), .B1(n1167), .Y(n41) );
  AOI31XL U584 ( .A0(n970), .A1(n971), .A2(n972), .B0(n911), .Y(n966) );
  AOI22XL U606 ( .A0(r2_out[2]), .A1(n914), .B0(n984), .B1(n1167), .Y(n107) );
  OAI21XL U747 ( .A0(top[3]), .A1(n951), .B0(n1066), .Y(n1063) );
  INVX1 U748 ( .A(newVal[4]), .Y(n1030) );
  NAND2X1 U749 ( .A(newVal[0]), .B(newVal[1]), .Y(n1012) );
  INVX1 U750 ( .A(newVal[1]), .Y(n1014) );
  INVX1 U751 ( .A(newVal[0]), .Y(n1013) );
  OAI21XL U752 ( .A0(r6_out[7]), .A1(n960), .B0(n1001), .Y(n1000) );
  OAI222XL U753 ( .A0(n960), .A1(r2_out[7]), .B0(n960), .B1(n1072), .C0(
        r2_out[7]), .C1(n1072), .Y(n997) );
  INVX1 U754 ( .A(n1073), .Y(n1072) );
  NOR2BX1 U755 ( .AN(r4_out[6]), .B(newVal[6]), .Y(n1045) );
  OAI21XL U756 ( .A0(newVal[4]), .A1(n1160), .B0(n1052), .Y(n1050) );
  NOR2BX1 U757 ( .AN(n991), .B(n998), .Y(n990) );
  AOI222X1 U758 ( .A0(newVal[7]), .A1(n1156), .B0(newVal[7]), .B1(n1059), .C0(
        n1156), .C1(n1059), .Y(n972) );
  OAI21XL U759 ( .A0(top[6]), .A1(n920), .B0(n1060), .Y(n1059) );
  OAI21XL U760 ( .A0(newVal[6]), .A1(n1161), .B0(n1061), .Y(n1060) );
  NOR2X1 U761 ( .A(n997), .B(n983), .Y(n991) );
  INVX1 U762 ( .A(n989), .Y(n979) );
  INVX1 U763 ( .A(clear), .Y(n993) );
  INVX1 U764 ( .A(n972), .Y(n983) );
  NAND2X1 U765 ( .A(n990), .B(n971), .Y(n996) );
  NAND2X1 U766 ( .A(n993), .B(n910), .Y(n981) );
  INVX1 U767 ( .A(newVal[2]), .Y(n987) );
  INVX1 U768 ( .A(newVal[3]), .Y(n951) );
  INVX1 U769 ( .A(n912), .Y(n935) );
  INVX1 U770 ( .A(newVal[5]), .Y(n937) );
  INVX1 U771 ( .A(newVal[7]), .Y(n960) );
  NAND2X1 U772 ( .A(loadIn), .B(n983), .Y(n918) );
  INVX1 U773 ( .A(newVal[6]), .Y(n920) );
  INVX1 U774 ( .A(n918), .Y(n940) );
  AOI21X1 U775 ( .A0(n1167), .A1(n980), .B0(clear), .Y(n914) );
  NOR2X1 U776 ( .A(n910), .B(n918), .Y(n924) );
  OAI21XL U777 ( .A0(n983), .A1(n969), .B0(n981), .Y(n922) );
  NOR2X1 U778 ( .A(loadIn), .B(n910), .Y(n923) );
  OAI21XL U779 ( .A0(n979), .A1(n911), .B0(n935), .Y(n927) );
  NOR2X1 U780 ( .A(n911), .B(n991), .Y(n912) );
  NOR2X1 U781 ( .A(n979), .B(n980), .Y(n913) );
  OAI21XL U782 ( .A0(n969), .A1(n927), .B0(n981), .Y(n908) );
  OAI21XL U783 ( .A0(n970), .A1(n995), .B0(n918), .Y(n931) );
  NOR3BX1 U784 ( .AN(n970), .B(n983), .C(n995), .Y(n932) );
  INVX1 U785 ( .A(loadIn), .Y(n911) );
  OAI21XL U786 ( .A0(n996), .A1(n969), .B0(n981), .Y(n929) );
  INVXL U787 ( .A(r5_out[4]), .Y(n1085) );
  OAI21XL U788 ( .A0(n1012), .A1(r5_out[0]), .B0(r5_out[1]), .Y(n1086) );
  OAI21XL U789 ( .A0(n1013), .A1(r5_out[0]), .B0(n1014), .Y(n1087) );
  NAND2X1 U790 ( .A(n951), .B(r5_out[3]), .Y(n1088) );
  NAND3X1 U791 ( .A(n1088), .B(n1086), .C(n1087), .Y(n1089) );
  AOI21X1 U792 ( .A0(n987), .A1(r5_out[2]), .B0(n1089), .Y(n1090) );
  OAI21XL U793 ( .A0(newVal[3]), .A1(n1159), .B0(newVal[2]), .Y(n1091) );
  OAI22X1 U794 ( .A0(r5_out[2]), .A1(n1091), .B0(r5_out[4]), .B1(n1030), .Y(
        n1092) );
  AOI211X1 U795 ( .A0(newVal[3]), .A1(n1159), .B0(n1090), .C0(n1092), .Y(n1093) );
  AOI21X1 U796 ( .A0(r5_out[5]), .A1(n937), .B0(n1093), .Y(n1094) );
  OAI21XL U797 ( .A0(newVal[4]), .A1(n1085), .B0(n1094), .Y(n1095) );
  OAI21XL U798 ( .A0(n937), .A1(r5_out[5]), .B0(n1095), .Y(n1096) );
  OAI2BB1X1 U799 ( .A0N(r5_out[6]), .A1N(n920), .B0(n1096), .Y(n1097) );
  OAI21XL U800 ( .A0(r5_out[6]), .A1(n920), .B0(n1097), .Y(n1098) );
  AOI222X1 U801 ( .A0(n1166), .A1(newVal[7]), .B0(n1166), .B1(n1098), .C0(
        newVal[7]), .C1(n1098), .Y(n971) );
  OAI21XL U802 ( .A0(newVal[3]), .A1(n1153), .B0(newVal[2]), .Y(n1099) );
  AOI222X1 U803 ( .A0(r2_out[2]), .A1(n1080), .B0(r2_out[2]), .B1(n987), .C0(
        n1080), .C1(n1099), .Y(n1079) );
  AOI21X1 U804 ( .A0(n1063), .A1(newVal[4]), .B0(n1065), .Y(n1100) );
  AOI222X1 U805 ( .A0(n937), .A1(top[5]), .B0(n937), .B1(n1100), .C0(top[5]), 
        .C1(n1100), .Y(n1061) );
  NAND2X1 U806 ( .A(r6_out[7]), .B(n960), .Y(n1101) );
  AOI21X1 U807 ( .A0(n1101), .A1(n1000), .B0(n996), .Y(n967) );
  AOI31X1 U808 ( .A0(n993), .A1(n990), .A2(loadIn), .B0(n968), .Y(n1102) );
  INVXL U809 ( .A(n1102), .Y(n925) );
  OAI21XL U810 ( .A0(newVal[5]), .A1(n1155), .B0(n1075), .Y(n1103) );
  AOI222X1 U811 ( .A0(r2_out[6]), .A1(n920), .B0(r2_out[6]), .B1(n1103), .C0(
        n920), .C1(n1103), .Y(n1073) );
  AOI22X1 U812 ( .A0(newVal[7]), .A1(n1165), .B0(n1157), .B1(newVal[6]), .Y(
        n1104) );
  OAI21XL U813 ( .A0(r3_out[3]), .A1(n951), .B0(n1039), .Y(n1105) );
  AOI2BB2X1 U814 ( .B0(newVal[4]), .B1(n1105), .A0N(n937), .A1N(r3_out[5]), 
        .Y(n1106) );
  INVXL U815 ( .A(r3_out[4]), .Y(n1107) );
  OAI21XL U816 ( .A0(newVal[4]), .A1(n1105), .B0(n1107), .Y(n1108) );
  AOI22X1 U817 ( .A0(n937), .A1(r3_out[5]), .B0(n1106), .B1(n1108), .Y(n1109)
         );
  OAI21XL U818 ( .A0(n1157), .A1(newVal[6]), .B0(n1109), .Y(n1110) );
  AOI22X1 U819 ( .A0(n960), .A1(r3_out[7]), .B0(n1104), .B1(n1110), .Y(n989)
         );
  AOI31X1 U820 ( .A0(n966), .A1(n967), .A2(n1167), .B0(n968), .Y(n1111) );
  INVXL U821 ( .A(n1111), .Y(n907) );
  INVXL U822 ( .A(newVal[3]), .Y(n1112) );
  OAI21XL U823 ( .A0(n1012), .A1(r3_out[0]), .B0(r3_out[1]), .Y(n1113) );
  NOR2X1 U824 ( .A(n1013), .B(r3_out[0]), .Y(n1114) );
  OAI21XL U825 ( .A0(n1114), .A1(newVal[1]), .B0(n1113), .Y(n1115) );
  AOI21X1 U826 ( .A0(r3_out[3]), .A1(n1112), .B0(n1115), .Y(n1116) );
  AOI21X1 U827 ( .A0(n951), .A1(r3_out[3]), .B0(n987), .Y(n1117) );
  AOI222X1 U828 ( .A0(n1163), .A1(n1116), .B0(n1163), .B1(n1117), .C0(n1116), 
        .C1(newVal[2]), .Y(n1039) );
  AND3X1 U829 ( .A(n970), .B(n972), .C(n971), .Y(n1118) );
  NOR3X1 U830 ( .A(n967), .B(n1118), .C(n969), .Y(n905) );
  INVX1 U831 ( .A(n910), .Y(n1167) );
  OAI21XL U832 ( .A0(loadIn), .A1(shiftOut), .B0(n993), .Y(n910) );
  INVX1 U833 ( .A(\r6/N1 ), .Y(n1168) );
endmodule

