library verilog;
use verilog.vl_types.all;
entity HEXtoSevenSeg is
    port(
        led             : out    vl_logic_vector(7 downto 0);
        digit           : in     vl_logic_vector(3 downto 0)
    );
end HEXtoSevenSeg;
