library verilog;
use verilog.vl_types.all;
entity finalTop is
end finalTop;
