library verilog;
use verilog.vl_types.all;
entity top1 is
end top1;
