library verilog;
use verilog.vl_types.all;
entity constants_sv_unit is
end constants_sv_unit;
