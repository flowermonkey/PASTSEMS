library verilog;
use verilog.vl_types.all;
entity toptest is
end toptest;
