library verilog;
use verilog.vl_types.all;
entity top_task3 is
end top_task3;
