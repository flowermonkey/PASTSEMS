library verilog;
use verilog.vl_types.all;
entity p18240_sv_unit is
end p18240_sv_unit;
